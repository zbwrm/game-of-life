`timescale 1ns / 1ps

module IS_3(
  input  Tl,T,Tr, L, R, Bl, B,Br, // Input Operands
  output Checked); 

  parameter DLY = 1;
  wire c1,c2,c3,c4,c5,c6,c7,c8,c9,c10;
  wire c11,c12,c13,c14,c15,c16,c17,c18;
  wire c19,c20,c21,c22,c23,c24,c25,c26;
  wire c27, c28,c29,c30,c31,c32,c33,c34;
  wire c35,c36,c37,c38,c39,c40,c41,c42,c43;
  wire c44, c45,c46,c47,c48,c49,c50,c51,c52;
  wire c53,c54,c55,c56;
  
  wire xor1, xor2, xor3, xor4, xor5;
  wire xor6, xor7, xor8, xor9, xor10;
  wire xor11, xor12, xor13, xor14, xor15;
  wire xor16, xor17, xor18, xor19, xor20;
  wire xor21, xor22, xor23, xor24, xor25;
  wire xor26, xor27, xor28, xor29, xor30;
  wire xor31, xor32, xor33, xor34, xor35;
  wire xor36, xor37, xor38, xor39, xor40;
  wire xor41, xor42, xor43, xor44, xor45;
  wire xor46, xor47, xor48, xor49, xor50;
  wire xor51, xor52, xor53, xor54;

  and #DLY G1(c1,Tl,T,Tr);
  and #DLY G2(c2,Tl,T,L);
  and #DLY G3(c3,Tl,T,R);
  and #DLY G4(c4,Tl,T,Bl);
  and #DLY G5(c5,Tl,T,B);
  and #DLY G6(c6,Tl,T,Br);
  and #DLY G7(c7,Tl,Tr,L);
  and #DLY G8(c8,Tl,Tr,R);
  and #DLY G9(c9,Tl,Tr,Bl);
  and #DLY G10(c10,Tl,Tr,B);
  and #DLY G11(c11,Tl,Tr,Br);
  and #DLY G12(c12,Tl,L,R);
  and #DLY G13(c13,Tl,L,Bl);
  and #DLY G14(c14,Tl,L,B);
  and #DLY G15(c15,Tl,L,Br);
  and #DLY G16(c16,Tl,R,Bl);
  and #DLY G17(c17,Tl,R,B);
  and #DLY G18(c18,Tl,R,Br);
  and #DLY G19(c19,Tl,Bl,B);
  and #DLY G20(c20,Tl,Bl,Br);
  and #DLY G21(c21,Tl,B,Br);
  and #DLY G22(c22,T,Tr,L);
  and #DLY G23(c23,T,Tr,R);
  and #DLY G24(c24,T,Tr,Bl);
  and #DLY G25(c25,T,Tr,B);
  and #DLY G26(c26,T,Tr,Br);
  and #DLY G27(c27,T,L,R);
  and #DLY G28(c28,T,L,Bl);
  and #DLY G29(c29,T,L,B);
  and #DLY G30(c30,T,L,Br);
  and #DLY G31(c31,T,R,Bl);
  and #DLY G32(c32,T,R,B);
  and #DLY G33(c33,T,R,Br);
  and #DLY G34(c34,T,Bl,B);
  and #DLY G35(c35,T,Bl,Br);
  and #DLY G36(c36,T,B,Br);
  and #DLY G37(c37,Tr,L,R);
  and #DLY G38(c38,Tr,L,Bl);
  and #DLY G39(c39,Tr,L,B);
  and #DLY G40(c40,Tr,L,Br);
  and #DLY G41(c41,Tr,R,Bl);
  and #DLY G42(c42,Tr,R,B);
  and #DLY G43(c43,Tr,R,Br);
  and #DLY G44(c44,Tr,Bl,B);
  and #DLY G45(c45,Tr,Bl,Br);
  and #DLY G46(c46,Tr,B,Br);
  and #DLY G47(c47,L,R,Bl);
  and #DLY G48(c48,L,R,B);
  and #DLY G49(c49,L,R,Br);
  and #DLY G50(c50,L,Bl,B);
  and #DLY G51(c51,L,Bl,Br);
  and #DLY G52(c52,L,B,Br);
  and #DLY G53(c53,R,Bl,B);
  and #DLY G54(c54,R,Bl,Br);
  and #DLY G55(c55,R,B,Br);
  and #DLY G56(c56,Bl,B,Br);
  
  xor #DLY xor_gate1(xor1, c1, c2);
  xor #DLY xor_gate2(xor2, c3, xor1);
  xor #DLY xor_gate3(xor3, c4, xor2);
  xor #DLY xor_gate4(xor4, c5, xor3);
  xor #DLY xor_gate5(xor5, c6, xor4);
  xor #DLY xor_gate6(xor6, c7, xor5);
  xor #DLY xor_gate7(xor7, c8, xor6);
  xor #DLY xor_gate8(xor8, c9, xor7);
  xor #DLY xor_gate9(xor9, c10, xor8);
  xor #DLY xor_gate10(xor10, c11, xor9);
  xor #DLY xor_gate11(xor11, c12, xor10);
  xor #DLY xor_gate12(xor12, c13, xor11);
  xor #DLY xor_gate13(xor13, c14, xor12);
  xor #DLY xor_gate14(xor14, c15, xor13);
  xor #DLY xor_gate15(xor15, c16, xor14);
  xor #DLY xor_gate16(xor16, c17, xor15);
  xor #DLY xor_gate17(xor17, c18, xor16);
  xor #DLY xor_gate18(xor18, c19, xor17);
  xor #DLY xor_gate19(xor19, c20, xor18);
  xor #DLY xor_gate20(xor20, c21, xor19);
  xor #DLY xor_gate21(xor21, c22, xor20);
  xor #DLY xor_gate22(xor22, c23, xor21);
  xor #DLY xor_gate23(xor23, c24, xor22);
  xor #DLY xor_gate24(xor24, c25, xor23);
  xor #DLY xor_gate25(xor25, c26, xor24);
  xor #DLY xor_gate26(xor26, c27, xor25);
  xor #DLY xor_gate27(xor27, c28, xor26);
  xor #DLY xor_gate28(xor28, c29, xor27);
  xor #DLY xor_gate29(xor29, c30, xor28);
  xor #DLY xor_gate30(xor30, c31, xor29);
  xor #DLY xor_gate31(xor31, c32, xor30);
  xor #DLY xor_gate32(xor32, c33, xor31);
  xor #DLY xor_gate33(xor33, c34, xor32);
  xor #DLY xor_gate34(xor34, c35, xor33);
  xor #DLY xor_gate35(xor35, c36, xor34);
  xor #DLY xor_gate36(xor36, c37, xor35);
  xor #DLY xor_gate37(xor37, c38, xor36);
  xor #DLY xor_gate38(xor38, c39, xor37);
  xor #DLY xor_gate39(xor39, c40, xor38);
  xor #DLY xor_gate40(xor40, c41, xor39);
  xor #DLY xor_gate41(xor41, c42, xor40);
  xor #DLY xor_gate42(xor42, c43, xor41);
  xor #DLY xor_gate43(xor43, c44, xor42);
  xor #DLY xor_gate44(xor44, c45, xor43);
  xor #DLY xor_gate45(xor45, c46, xor44);
  xor #DLY xor_gate46(xor46, c47, xor45);
  xor #DLY xor_gate47(xor47, c48, xor46);
  xor #DLY xor_gate48(xor48, c49, xor47);
  xor #DLY xor_gate49(xor49, c50, xor48);
  xor #DLY xor_gate50(xor50, c51, xor49);
  xor #DLY xor_gate51(xor51, c52, xor50);
  xor #DLY xor_gate52(xor52, c53, xor51);
  xor #DLY xor_gate53(xor53, c54, xor52);
  xor #DLY xor_gate54(xor54, c55, xor53);
  xor #DLY xor_gate55(Checked, c56, xor54);
endmodule
